module Snooping (clock);

maquinaSnooping maquina();	

endmodule
