module Tomasulo (Clock);

	input Clock;
	
	controle_RS control (Clock);

endmodule
