module testeMaquina ();

maquinaUnica maquina(maquina, op, estadoAtual, entradaBarramento, novoEstado, saidaBarramento, writeBack, abortAccessMemory);